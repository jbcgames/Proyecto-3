// **********************
// Multiplier Unit Module
// **********************
module multiplierunit (dataA, dataB, dataR);
	input logic [31:0] dataA, dataB;
	output logic [31:0] dataR;

	// Internal signals to perform the multiplication
	// WRITE HERE YOUR CODE
			
	// Process: sign XORer
	// WRITE HERE YOUR CODE
	
	// Process: exponent adder
	// WRITE HERE YOUR CODE
	
	// Process: mantissa multiplier
	// WRITE HERE YOUR CODE
	
	// Process: operand validator and result normalizer and assembler
	// WRITE HERE YOUR CODE
endmodule

// ***************************** 
// Testbench for Multiplier Unit
// ***************************** 
module tb_multiplierunit ();
	// WRITE HERE YOUR CODE
endmodule