// *******************
// Control Unit Module
// *******************
module controlunit (clk, rst, loaddata, inputdata_ready, boton, led);
	input logic  clk, rst, boton;
	output logic  loaddata;
	output logic [3:0]led;
	input logic inputdata_ready;
	logic senal, reset;
	pulse Pulso(clk, rst, boton, senal);
	typedef enum logic [3:0] {A1, A2, A3, A4, B1, B2, B3, B4, R1, R2, R3, R4} State;
	State momento;
	always_comb begin
	reset=~rst;
	end
	always_ff @(posedge reset, posedge senal)begin
	if(reset)begin
	momento<=A1;
	end else if(momento==A1)begin
	momento<=A2;
	end else if(momento==A2)begin
	momento<=A3;
	end else if(momento==A3)begin
	momento<=A4;
	end else if(momento==A4)begin
	momento<=B1;
	end else if(momento==B1)begin
	momento<=B2;
	end else if(momento==B2)begin
	momento<=B3;
	end else if(momento==B3)begin
	momento<=B4;
	end else if(momento==B4)begin
	momento<=R1;
	end else if(momento==R1)begin
	momento<=R2;
	end else if(momento==R2)begin
	momento<=R3;
	end else if(momento==R3)begin
	momento<=R4;
	end else if(momento==R4)begin
	momento<=R1;
	end
	end
	
 always_comb begin
 case(momento)
	 A1:led=4'b0001;
	 A2:led=4'b0010;
	 A3:led=4'b0011;
	 A4:led=4'b0100;
	 B1:led=4'b0101;
	 B2:led=4'b0110;
	 B3:led=4'b0111;
	 B4:led=4'b1000;
	 R1:led=4'b1001;
	 R2:led=4'b1010;
	 R3:led=4'b1011;
	 R4:led=4'b1100;
endcase
 end
 
endmodule

